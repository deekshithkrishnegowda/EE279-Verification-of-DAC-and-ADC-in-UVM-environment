//package test_package ;

//import uvm_pkg ::*;

`include "uvm_macros.svh"

//`include "../top/dut_intf.sv"
`include "../uvo/messages.sv"
`include "../uvo/sequence.sv"
`include "../uvc/driver.sv"
`include "../uvc/sequencer.sv"
`include "../uvc/monitor_dac0.sv"
`include "../uvc/monitor_dac1.sv"

`include "../uvc/bfm.sv"
`include "../uvc/monitor_adc0.sv"
`include "../uvc/monitor_adc1.sv"

`include "../uvc/agent.sv"
`include "../uvc/virtual_sequencer.sv"
`include "../uvc/virtual_sequence.sv"
`include "../uvc/scoreboard.sv"
`include "../uvc/environment.sv"
`include "../uvc/test.sv"



//endpackage
